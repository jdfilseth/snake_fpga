/*
Based off the VGA controller file in DE-10 lite demonstration, but heavily modified for snake game
*/

module vga_controller(vga_reset,
                      vga_clk,
					  board_state,
					  is_start_screen,
					  is_over,
                      oHS,
                      oVS,
                      oVGA_B,
                      oVGA_G,
                      oVGA_R);
					  
`include "game_vga_param.h"	  


			
input vga_reset;
input vga_clk;
input is_start_screen;
input is_over;
input [39*29*3-1:0] board_state;

output reg oHS;
output reg oVS;
output [3:0] oVGA_B;
output [3:0] oVGA_G;  
output [3:0] oVGA_R;                       
///////// ////                     
reg [18:0] h_addr ;
reg [18:0] v_addr ;
reg inc_vert;
wire [7:0] index;
wire [23:0] bgr_data_raw;
wire cBLANK_n,cVBLANK_n,cHS,cVS,rst;
////
assign rst = ~vga_reset;

reg [11:0] bgr_data;

wire [BOARD_HEIGHT_BITS-1:0] v_cell;
wire [BOARD_WIDTH_BITS-1:0] h_cell;
wire [3:0] v_pos, h_pos;
wire [8:0] sq_dist_from_ctr;

// locations of cells in screen, and individual units within cells
assign v_cell = (v_addr + 8)/CELL_SIZE;
assign h_cell = (h_addr + 8)/CELL_SIZE;
assign v_pos = (v_addr + 8)%CELL_SIZE;
assign h_pos = (h_addr + 8)%CELL_SIZE;
assign sq_dist_from_ctr = (v_pos-8)*(v_pos-8) + (h_pos-8)*(h_pos-8);

// restructure board state into more easily usable array format
wire[3:0] board_state_wires [BOARD_WIDTH:1][BOARD_HEIGHT:1];

genvar v;
generate 
	for (v=0; v<29*39; v=v+1) begin : boardgen
		assign board_state_wires[v/29 + 1][v%29 + 1] = board_state[v*3+2:v*3];
	end
endgenerate


wire [0:START_SCREEN_W*START_SCREEN_H-1] start_screen;
wire [0:GAME_OVER_ARR_W*GAME_OVER_ARR_H-1] game_over_screen;



video_sync_generator LTM_ins (.vga_clk(vga_clk),
                              .reset(rst),
                              .blank_n(cBLANK_n),
							  .vblank_n(cVBLANK_n),
                              .HS(cHS),
                              .VS(cVS)
										);

////Address generator
always@(posedge vga_clk,negedge vga_reset)
begin
  if (!vga_reset)
  begin
     h_addr<=19'd0;
	 v_addr<=19'd0;
	 inc_vert<=1;
  end
  else 
  begin
	if (cBLANK_n==1'b1)
	begin
		h_addr<=h_addr+1;
		inc_vert<=1;
	end
	else
	begin
		h_addr<=19'd0;
		if (cVBLANK_n==1'b1)
		begin
			if (inc_vert==1)
			begin
				v_addr<=v_addr+1;
				inc_vert<=0;
			end
		end
		else
			v_addr<=19'd0;
	end

  end
  

  
end

// VGA output colors
always@(posedge vga_clk)
begin
	if (~vga_reset)
    	bgr_data<=12'h000;
	
	// draw gray border at edge of monitor
    else if (v_cell==0 || v_cell==BOARD_HEIGHT+1 || h_cell==0 || h_cell==BOARD_WIDTH+1)
		bgr_data <= {4'hc, 4'hc, 4'hc};
		
	// main game board
	else if (v_cell > 0 && v_cell < BOARD_HEIGHT+1 && h_cell > 0 && h_cell < BOARD_WIDTH+1)
	begin
		// draw start screen
		if (is_start_screen)
		begin
			if (
				(h_addr < (VIDEO_W - START_SCREEN_W)/2 - MESSAGE_BORDER) || (h_addr >= (START_SCREEN_W + VIDEO_W)/2 + MESSAGE_BORDER) ||
				(v_addr < (VIDEO_H - START_SCREEN_H)/2 - MESSAGE_BORDER) || (v_addr >= (START_SCREEN_H + VIDEO_H)/2 + MESSAGE_BORDER)
			)
				bgr_data <= 12'h000;
			else if (
				(h_addr < (VIDEO_W - START_SCREEN_W)/2) || (h_addr >= (START_SCREEN_W + VIDEO_W)/2) ||
				(v_addr < (VIDEO_H - START_SCREEN_H)/2) || (v_addr >= (START_SCREEN_H + VIDEO_H)/2)
			)
				bgr_data <= 12'hf00;
			else if (start_screen[(v_addr - (VIDEO_H - START_SCREEN_H)/2)*START_SCREEN_W + h_addr - (VIDEO_W - START_SCREEN_W)/2]==1)
				bgr_data <= 12'h00f;
			else
				bgr_data <= 12'hf00;			
		end
		
		// draw game over screen on top of game
		else if (is_over && 
			!(
				(h_addr < (VIDEO_W - GAME_OVER_ARR_W)/2 - MESSAGE_BORDER) || (h_addr >= (GAME_OVER_ARR_W + VIDEO_W)/2 + MESSAGE_BORDER) ||
				(v_addr < (VIDEO_H - GAME_OVER_ARR_H)/2 - MESSAGE_BORDER) || (v_addr >= (GAME_OVER_ARR_H + VIDEO_H)/2 + MESSAGE_BORDER)
			)
		)
		begin
			if (
				(h_addr < (VIDEO_W - GAME_OVER_ARR_W)/2) || (h_addr >= (GAME_OVER_ARR_W + VIDEO_W)/2) ||
				(v_addr < (VIDEO_H - GAME_OVER_ARR_H)/2) || (v_addr >= (GAME_OVER_ARR_H + VIDEO_H)/2)
			)
				bgr_data <= 12'hf00;
			else if (game_over_screen[(v_addr - (VIDEO_H - GAME_OVER_ARR_H)/2)*GAME_OVER_ARR_W + h_addr - (VIDEO_W - GAME_OVER_ARR_W)/2]==1)
				bgr_data <= 12'h00f;
			else
				bgr_data <= 12'hf00;			
		end
		
		// draw rest of board based on board_state_wires
		else
		begin
			// draw black border around snake segments
			if (v_pos < 1 || v_pos >= 15 || h_pos < 1 || h_pos >= 15)
				bgr_data <= 12'h000;
			else
			begin
				// draw green snake segments
				if (board_state_wires[h_cell][v_cell]>0 && board_state_wires[h_cell][v_cell]<7)
					bgr_data <= 12'h0f0;

				else if (board_state_wires[h_cell][v_cell]==7)
				begin
					
					// draw yellow dots
					if (sq_dist_from_ctr < 25)
						bgr_data <= 12'h0ff;

					else
						bgr_data <= 12'h000;
				end
				else
					bgr_data <= 12'h000;
			end
		end
	end
	else
		bgr_data <= 12'h000; 
end

assign oVGA_B=bgr_data[11:8];
assign oVGA_G=bgr_data[7:4]; 
assign oVGA_R=bgr_data[3:0];
///////////////////
//////Delay the iHD, iVD,iDEN for one clock cycle;
reg mHS, mVS;
always@(posedge vga_clk)
begin
  mHS<=cHS;
  mVS<=cVS;
  oHS<=mHS;
  oVS<=mVS;
end

// parameters need to match dimensions of arrays below
parameter   START_SCREEN_W 		= 315;
parameter	START_SCREEN_H 		= 97;
parameter	GAME_OVER_ARR_W 	= 354;
parameter	GAME_OVER_ARR_H 	= 96;

// start screen message
assign start_screen = {
315'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111000000000000000000000000011111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000,
315'b000000000000000000000000000000000111111000000000000001111110000000000000111111000111111111111111111111111000011111100000000000000000000000000111111111111110000000000000000111111111111100000000000000011111111000000000000000001111111000000111111111111111111111111000000011111000000000000000000000000000000000000000000,
315'b000000000000000000000000000000000011111000000000000001111110000000000000111111000111111111111111111111111000011111100000000000000000000000001111111111111111110000000000011111111111111111000000000000011111111000000000000000011111111000000111111111111111111111111000000011111000000000000000000000000000000000000000000,
315'b000000000000000000000000000000000011111000000000000011111110000000000000111110000111111111111111111111111000011111100000000000000000000000111111111111111111111000000000111111111111111111110000000000011111111100000000000000011111111000000111111111111111111111111000000011111000000000000000000000000000000000000000000,
315'b000000000000000000000000000000000011111100000000000011111110000000000000111110000111111111111111111111111000011111100000000000000000000001111111111111111111111100000011111111111111111111111000000000011111111100000000000000111111111000000111111111111111111111111000000011111000000000000000000000000000000000000000000,
315'b000000000000000000000000000000000011111100000000000011111111000000000001111110000111111111111111111111111000011111100000000000000000000011111111100000011111111100000111111111100000011111111100000000011111111110000000000000111111111000000111111111111111111111111000000011111000000000000000000000000000000000000000000,
315'b000000000000000000000000000000000001111100000000000011111111000000000001111110000111111000000000000000000000011111100000000000000000000111111110000000000011111100000111111110000000000111111110000000011111111110000000000001111111111000000111111000000000000000000000000011111000000000000000000000000000000000000000000,
315'b000000000000000000000000000000000001111100000000000111111111000000000001111100000111111000000000000000000000011111100000000000000000001111111100000000000000111100001111111000000000000011111110000000011111111110000000000001111111111000000111111000000000000000000000000011111000000000000000000000000000000000000000000,
315'b000000000000000000000000000000000001111110000000000111111111000000000001111100000111111000000000000000000000011111100000000000000000001111111000000000000000011100001111110000000000000001111111000000011111111111000000000001111111111000000111111000000000000000000000000011111000000000000000000000000000000000000000000,
315'b000000000000000000000000000000000001111110000000000111111111000000000011111100000111111000000000000000000000011111100000000000000000011111110000000000000000001000011111100000000000000000111111000000011111111111000000000011111011111000000111111000000000000000000000000011111000000000000000000000000000000000000000000,
315'b000000000000000000000000000000000000111110000000000111101111100000000011111100000111111000000000000000000000011111100000000000000000011111100000000000000000000000011111100000000000000000011111100000011111101111100000000011111011111000000111111000000000000000000000000011111000000000000000000000000000000000000000000,
315'b000000000000000000000000000000000000111110000000001111101111100000000011111000000111111000000000000000000000011111100000000000000000111111100000000000000000000000111111000000000000000000011111100000011111101111100000000111110011111000000111111000000000000000000000000011111000000000000000000000000000000000000000000,
315'b000000000000000000000000000000000000111111000000001111101111100000000011111000000111111000000000000000000000011111100000000000000000111111000000000000000000000000111111000000000000000000011111100000011111100111110000000111110011111000000111111000000000000000000000000011111000000000000000000000000000000000000000000,
315'b000000000000000000000000000000000000111111000000001111000111100000000011111000000111111000000000000000000000011111100000000000000000111111000000000000000000000000111111000000000000000000001111100000011111100111110000001111100011111000000111111000000000000000000000000011111000000000000000000000000000000000000000000,
315'b000000000000000000000000000000000000011111000000001111000111110000000111111000000111111000000000000000000000011111100000000000000000111111000000000000000000000000111111000000000000000000001111110000011111100111111000001111100011111000000111111000000000000000000000000011111000000000000000000000000000000000000000000,
315'b000000000000000000000000000000000000011111000000011111000111110000000111110000000111111111111111111111110000011111100000000000000000111110000000000000000000000000111110000000000000000000001111110000011111100011111000001111000011111000000111111111111111111111110000000011111000000000000000000000000000000000000000000,
315'b000000000000000000000000000000000000011111100000011111000111110000000111110000000111111111111111111111110000011111100000000000000000111110000000000000000000000001111110000000000000000000001111110000011111100011111100011111000011111000000111111111111111111111110000000011111000000000000000000000000000000000000000000,
315'b000000000000000000000000000000000000011111100000011110000011110000000111110000000111111111111111111111110000011111100000000000000001111110000000000000000000000001111110000000000000000000001111110000011111100001111100011111000011111000000111111111111111111111110000000011111000000000000000000000000000000000000000000,
315'b000000000000000000000000000000000000001111100000011110000011111000001111110000000111111111111111111111110000011111100000000000000001111110000000000000000000000001111110000000000000000000001111110000011111100001111100111110000011111000000111111111111111111111110000000011111000000000000000000000000000000000000000000,
315'b000000000000000000000000000000000000001111100000111110000011111000001111100000000111111111111111111111110000011111100000000000000001111110000000000000000000000001111110000000000000000000001111110000011111100000111110111110000011111000000111111111111111111111110000000011111000000000000000000000000000000000000000000,
315'b000000000000000000000000000000000000001111110000111110000011111000001111100000000111111000000000000000000000011111100000000000000001111110000000000000000000000001111110000000000000000000001111110000011111100000111111111100000011111000000111111000000000000000000000000011111000000000000000000000000000000000000000000,
315'b000000000000000000000000000000000000001111110000111110000001111000001111100000000111111000000000000000000000011111100000000000000001111110000000000000000000000001111110000000000000000000001111110000011111100000111111111100000011111000000111111000000000000000000000000011111000000000000000000000000000000000000000000,
315'b000000000000000000000000000000000000000111110000111100000001111100011111100000000111111000000000000000000000011111100000000000000000111110000000000000000000000001111110000000000000000000001111110000011111100000011111111000000011111000000111111000000000000000000000000011111000000000000000000000000000000000000000000,
315'b000000000000000000000000000000000000000111110000111100000001111100011111000000000111111000000000000000000000011111100000000000000000111110000000000000000000000000111110000000000000000000001111110000011111100000011111111000000011111000000111111000000000000000000000000011111000000000000000000000000000000000000000000,
315'b000000000000000000000000000000000000000111111001111100000001111100011111000000000111111000000000000000000000011111100000000000000000111111000000000000000000000000111110000000000000000000001111110000011111100000001111110000000011111000000111111000000000000000000000000011111000000000000000000000000000000000000000000,
315'b000000000000000000000000000000000000000111111001111100000000111100011111000000000111111000000000000000000000011111100000000000000000111111000000000000000000000000111111000000000000000000001111100000011111100000001111110000000011111000000111111000000000000000000000000011111000000000000000000000000000000000000000000,
315'b000000000000000000000000000000000000000011111001111000000000111110111111000000000111111000000000000000000000011111100000000000000000111111000000000000000000000000111111000000000000000000011111100000011111100000000111110000000011111000000111111000000000000000000000000011111000000000000000000000000000000000000000000,
315'b000000000000000000000000000000000000000011111001111000000000111110111110000000000111111000000000000000000000011111100000000000000000111111100000000000000000000000111111000000000000000000011111100000011111100000000111100000000011111000000111111000000000000000000000000011111000000000000000000000000000000000000000000,
315'b000000000000000000000000000000000000000011111111111000000000111110111110000000000111111000000000000000000000011111100000000000000000011111100000000000000000000000011111100000000000000000011111100000011111100000000000000000000011111000000111111000000000000000000000000000000000000000000000000000000000000000000000000,
315'b000000000000000000000000000000000000000011111111111000000000011111111110000000000111111000000000000000000000011111100000000000000000011111110000000000000000001000011111110000000000000000111111000000011111100000000000000000000011111000000111111000000000000000000000000000000000000000000000000000000000000000000000000,
315'b000000000000000000000000000000000000000001111111110000000000011111111110000000000111111000000000000000000000011111100000000000000000001111111000000000000000011100001111110000000000000001111111000000011111100000000000000000000011111000000111111000000000000000000000000000000000000000000000000000000000000000000000000,
315'b000000000000000000000000000000000000000001111111110000000000011111111100000000000111111000000000000000000000011111100000000000000000001111111100000000000000111100001111111000000000000011111110000000011111100000000000000000000011111000000111111000000000000000000000000000000000000000000000000000000000000000000000000,
315'b000000000000000000000000000000000000000001111111110000000000011111111100000000000111111000000000000000000000011111100000000000000000000111111110000000000011111100000111111110000000000111111110000000011111100000000000000000000011111000000111111000000000000000000000000011111000000000000000000000000000000000000000000,
315'b000000000000000000000000000000000000000000111111110000000000001111111100000000000111111111111111111111111000011111111111111111111110000011111111100000011111111100000111111111100000011111111100000000011111100000000000000000000011111000000111111111111111111111111000000011111000000000000000000000000000000000000000000,
315'b000000000000000000000000000000000000000000111111100000000000001111111100000000000111111111111111111111111000011111111111111111111110000001111111111111111111111100000011111111111111111111111000000000011111100000000000000000000011111000000111111111111111111111111000000011111000000000000000000000000000000000000000000,
315'b000000000000000000000000000000000000000000111111100000000000001111111000000000000111111111111111111111111000011111111111111111111110000000111111111111111111111000000000111111111111111111110000000000011111100000000000000000000011111000000111111111111111111111111000000011111000000000000000000000000000000000000000000,
315'b000000000000000000000000000000000000000000111111100000000000001111111000000000000111111111111111111111111000011111111111111111111110000000011111111111111111100000000000011111111111111111000000000000011111100000000000000000000011111000000111111111111111111111111000000011111000000000000000000000000000000000000000000,
315'b000000000000000000000000000000000000000000011111100000000000000111111000000000000111111111111111111111111000011111111111111111111110000000000111111111111110000000000000000111111111111110000000000000011111000000000000000000000011111000000111111111111111111111111000000011111000000000000000000000000000000000000000000,
315'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111100000000000000000000000111111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000,
315'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000,
315'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000,
315'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000,
315'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000,
315'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000,
315'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000,
315'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000,
315'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000,
315'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000,
315'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000,
315'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000,
315'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000,
315'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000,
315'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000,
315'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000,
315'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000,
315'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000,
315'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000,
315'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000,
315'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000,
315'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000,
315'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000,
315'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000,
315'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000,
315'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000,
315'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000,
315'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000,
315'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000,
315'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000,
315'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000,
315'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000,
315'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000,
315'b111111111110000000011111111111000000000001111111111111111100000011111111110000000001111111111000000000000000001111000000000011110000000001110000000000000000000111111111111111111110000000111111111000000000000000000000000011111111110001111111111111111111100000001111100000000001111111111100000000111111111111111111110,
315'b111111111111100000011111111111111000000001111111111111111100001111111111111100000111111111111110000000000000001111000000000111110000000011110000000000000000000111111111111111111110000011111111111110000000000000000000001111111111111101111111111111111111100000001111100000000001111111111111100000111111111111111111110,
315'b111111111111111000011111111111111100000001111111111111111100011111111111111100001111111111111110000000000000001111000000001111100000000111110000000000000000000111111111111111111110000111111111111111000000000000000000011111111111111101111111111111111111100000011111110000000001111111111111110000111111111111111111110,
315'b111111111111111000011111111111111110000001111111111111111100111111000001111100011111100000111110000000000000001111000000011111000000011111110000000000000000000111111111111111111110001111110000011111100000000000000000111111000001111101111111111111111111100000011111110000000001111111111111111000111111111111111111110,
315'b111100000001111100011110000000111110000001111000000000000000111100000000011100011110000000001110000000000000001111000000111110000000111111110000000000000000000000000001111000000000011111000000000111110000000000000000111100000000011100000000011110000000000000011111110000000001111000000011111000000000001111000000000,
315'b111100000000111110011110000000011110000001111000000000000000111100000000000100011110000000000010000000000000001111000001111100000000111111110000000000000000000000000001111000000000011110000000000011110000000000000000111100000000000100000000011110000000000000111101111000000001111000000001111000000000001111000000000,
315'b111100000000011110011110000000001111000001111000000000000001111000000000000000111100000000000000000000000000001111000001111000000000000011110000000000000000000000000001111000000000111100000000000011111000000000000001111000000000000000000000011110000000000000111101111000000001111000000000111100000000001111000000000,
315'b111100000000011110011110000000001111000001111000000000000001111000000000000000111100000000000000000000000000001111000011110000000000000011110000000000000000000000000001111000000000111100000000000001111000000000000001111000000000000000000000011110000000000000111001111000000001111000000000111100000000001111000000000,
315'b111100000000011110011110000000001111000001111000000000000001111100000000000000111110000000000000000000000000001111000111100000000000000011110000000000000000000000000001111000000000111100000000000001111000000000000001111100000000000000000000011110000000000001111000111100000001111000000000111100000000001111000000000,
315'b111100000000011110011110000000011110000001111000000000000000111110000000000000011111000000000000000000000000001111001111000000000000000011110000000000000000000000000001111000000001111000000000000001111100000000000000111110000000000000000000011110000000000001111000111100000001111000000001111000000000001111000000000,
315'b111100000000111100011110000000011110000001111111111111111000111111100000000000011111110000000000000000000000001111011110000000000000000011110000000000000000000000000001111000000001111000000000000000111100000000000000111111100000000000000000011110000000000001111000111100000001111000000001111000000000001111000000000,
315'b111100000000111100011110000000111110000001111111111111111000011111111100000000001111111110000000000000000000001111111110000000000000000011110000000000000000000000000001111000000001111000000000000000111100000000000000011111111100000000000000011110000000000011110000011110000001111000000011111000000000001111000000000,
315'b111100000011111100011110000111111100000001111111111111111000001111111111100000000111111111110000000000000000001111111110000000000000000011110000000000000000000000000001111000000001111000000000000000111100000000000000001111111111100000000000011110000000000011110000011110000001111000011111110000000000001111000000000,
315'b111111111111111000011111111111111000000001111111111111111000000111111111111000000011111111111100000000000000001111111111000000000000000011110000000000000000000000000001111000000001111000000000000000111100000000000000000111111111111000000000011110000000000011110000011110000001111111111111100000000000001111000000000,
315'b111111111111110000011111111111100000000001111000000000000000000000111111111100000000011111111110000000000000001111111111100000000000000011110000000000000000000000000001111000000001111000000000000000111100000000000000000000111111111100000000011110000000000111100000001111000001111111111110000000000000001111000000000,
315'b111111111111000000011111111111100000000001111000000000000000000000000011111100000000000001111110000000000000001111001111100000000000000011110000000000000000000000000001111000000001111000000000000000111100000000000000000000000011111100000000011110000000000111100000001111000001111111111110000000000000001111000000000,
315'b111111100000000000011110000111110000000001111000000000000000000000000000111110000000000000011111000000000000001111000111110000000000000011110000000000000000000000000001111000000001111000000000000000111000000000000000000000000000111110000000011110000000000111111111111111000001111000011111000000000000001111000000000,
315'b111100000000000000011110000011111000000001111000000000000000000000000000111110000000000000011111000000000000001111000011111000000000000011110000000000000000000000000001111000000000111100000000000001111000000000000000000000000000111110000000011110000000001111111111111111100001111000001111100000000000001111000000000,
315'b111100000000000000011110000001111100000001111000000000000000000000000000011110000000000000001111000000000000001111000001111100000000000011110000000000000000000000000001111000000000111100000000000001111000000000000000000000000000011110000000011110000000001111111111111111100001111000000111110000000000001111000000000,
315'b111100000000000000011110000000111110000001111000000000000000000000000000011110000000000000001111000000000000001111000001111110000000000011110000000000000000000000000001111000000000111100000000000011111000000000000000000000000000011110000000011110000000001111000000000111100001111000000011111000000000001111000000000,
315'b111100000000000000011110000000111110000001111000000000000001100000000000011100110000000000001110000000000000001111000000111110000000000011110000000000000000000000000001111000000000011110000000000011110000000000000001100000000000011100000000011110000000011110000000000011110001111000000011111000000000001111000000000,
315'b111100000000000000011110000000011111000001111000000000000001110000000000111100111000000000011110000000000000001111000000011111000000000011110000000000000000000000000001111000000000011111000000000111110000000000000001110000000000111100000000011110000000011110000000000011110001111000000001111100000000001111000000000,
315'b111100000000000000011110000000001111100001111000000000000001111100000011111100111110000001111110000000000000001111000000001111100000000011110000000000000000000000000001111000000000001111110000011111100000000000000001111100000011111100000000011110000000011110000000000011110001111000000000111110000000001111000000000,
315'b111100000000000000011110000000000111110001111111111111111101111111111111111000111111111111111100000000000000001111000000000111110000111111111111000000000000000000000001111000000000001111111111111111000000000000000001111111111111111000000000011110000000111100000000000001111001111000000000011111000000001111000000000,
315'b111100000000000000011110000000000011111001111111111111111101111111111111110000111111111111111000000000000000001111000000000111110000111111111111000000000000000000000001111000000000000011111111111110000000000000000001111111111111110000000000011110000000111100000000000001111001111000000000001111100000001111000000000,
315'b111100000000000000011110000000000011111001111111111111111100001111111111000000000111111111100000000000000000001111000000000011111000111111111111000000000000000000000001111000000000000001111111111100000000000000000000001111111111000000000000011110000000111100000000000001111001111000000000001111100000001111000000000
};


assign game_over_screen = {
354'b000000000000000000000000000000000000000000000001111111111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111111111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000,
354'b000000000000000000000000000000000000000000001111111111111111000000000000000000111111000000000000000011111110000000000000000011111110000000111111111111111111111110000000000000000000000000000111111111111111000000000011111000000000000000000011111000011111111111111111111111000001111111111111111100000000000000001111100000000000000000000000000000000000000000,
354'b000000000000000000000000000000000000000000111111111111111111111000000000000001111111100000000000000011111110000000000000000111111110000000111111111111111111111110000000000000000000000000011111111111111111100000000011111000000000000000000011111000011111111111111111111111000001111111111111111111000000000000001111100000000000000000000000000000000000000000,
354'b000000000000000000000000000000000000000001111111111111111111111100000000000001111111100000000000000011111111000000000000000111111110000000111111111111111111111110000000000000000000000000111111111111111111111000000011111000000000000000000011110000011111111111111111111111000001111111111111111111100000000000001111100000000000000000000000000000000000000000,
354'b000000000000000000000000000000000000000011111111000000011111111100000000000001111111100000000000000011111111000000000000001111111110000000111111111111111111111110000000000000000000000001111111100000001111111100000001111100000000000000000111110000011111111111111111111111000001111111111111111111110000000000001111100000000000000000000000000000000000000000,
354'b000000000000000000000000000000000000000111111100000000000011111100000000000011111111110000000000000011111111100000000000001111111110000000111110000000000000000000000000000000000000000011111110000000000011111110000001111100000000000000000111110000011111000000000000000000000001111100000000001111111000000000001111100000000000000000000000000000000000000000,
354'b000000000000000000000000000000000000001111110000000000000000111100000000000011111111110000000000000011111111100000000000001111111110000000111110000000000000000000000000000000000000000111111000000000000001111110000001111100000000000000000111100000011111000000000000000000000001111100000000000111111000000000001111100000000000000000000000000000000000000000,
354'b000000000000000000000000000000000000011111100000000000000000001100000000000011110011110000000000000011110111100000000000011110111110000000111110000000000000000000000000000000000000000111110000000000000000111111000000111110000000000000001111100000011111000000000000000000000001111100000000000011111100000000001111100000000000000000000000000000000000000000,
354'b000000000000000000000000000000000000011111100000000000000000000100000000000111110011111000000000000011110011110000000000011110111110000000111110000000000000000000000000000000000000001111110000000000000000011111000000111110000000000000001111100000011111000000000000000000000001111100000000000001111100000000001111100000000000000000000000000000000000000000,
354'b000000000000000000000000000000000000111111000000000000000000000000000000000111110011111000000000000011110011110000000000111100111110000000111110000000000000000000000000000000000000001111100000000000000000011111100000111110000000000000001111000000011111000000000000000000000001111100000000000001111100000000001111100000000000000000000000000000000000000000,
354'b000000000000000000000000000000000000111110000000000000000000000000000000000111100001111000000000000011110011111000000000111100111110000000111110000000000000000000000000000000000000011111100000000000000000001111100000011111000000000000011111000000011111000000000000000000000001111100000000000001111100000000001111100000000000000000000000000000000000000000,
354'b000000000000000000000000000000000000111110000000000000000000000000000000001111100001111100000000000011110001111000000001111000111110000000111110000000000000000000000000000000000000011111000000000000000000001111100000011111000000000000011111000000011111000000000000000000000001111100000000000001111100000000001111100000000000000000000000000000000000000000,
354'b000000000000000000000000000000000001111100000000000000000000000000000000001111100001111100000000000011110001111100000001111000111110000000111110000000000000000000000000000000000000011111000000000000000000001111110000011111000000000000011110000000011111000000000000000000000001111100000000000001111100000000001111100000000000000000000000000000000000000000,
354'b000000000000000000000000000000000001111100000000000000000000000000000000001111000000111100000000000011110000111100000011110000111110000000111110000000000000000000000000000000000000011111000000000000000000000111110000001111100000000000111110000000011111000000000000000000000001111100000000000001111100000000001111100000000000000000000000000000000000000000,
354'b000000000000000000000000000000000001111100000000000000000000000000000000011111000000111110000000000011110000111110000011110000111110000000111110000000000000000000000000000000000000111110000000000000000000000111110000001111100000000000111110000000011111000000000000000000000001111100000000000011111000000000001111100000000000000000000000000000000000000000,
354'b000000000000000000000000000000000001111100000000000000000000000000000000011111000000111110000000000011110000011110000011110000111110000000111111111111111111111100000000000000000000111110000000000000000000000111110000001111100000000000111100000000011111111111111111111110000001111100000000000011111000000000001111100000000000000000000000000000000000000000,
354'b000000000000000000000000000000000001111100000000000000000000000000000000011110000000111110000000000011110000011110000111100000111110000000111111111111111111111100000000000000000000111110000000000000000000000111110000000111110000000001111100000000011111111111111111111110000001111100000000000111110000000000001111100000000000000000000000000000000000000000,
354'b000000000000000000000000000000000001111100000000000000000000000000000000111110000000011111000000000011110000011111000111100000111110000000111111111111111111111100000000000000000000111110000000000000000000000111110000000111110000000001111100000000011111111111111111111110000001111100000000011111110000000000001111100000000000000000000000000000000000000000,
354'b000000000000000000000000000000000001111100000000000000000000000000000000111110000000011111000000000011110000001111001111000000111110000000111111111111111111111100000000000000000000111110000000000000000000000111110000000111110000000001111000000000011111111111111111111110000001111111111111111111100000000000001111100000000000000000000000000000000000000000,
354'b000000000000000000000000000000000001111100000000000111111111111100000000111100000000011111000000000011110000001111101111000000111110000000111110000000000000000000000000000000000000111110000000000000000000000111110000000011111000000011111000000000011111000000000000000000000001111111111111111110000000000000001111100000000000000000000000000000000000000000,
354'b000000000000000000000000000000000001111100000000000111111111111100000001111100000000001111100000000011110000000111111110000000111110000000111110000000000000000000000000000000000000111110000000000000000000000111110000000011111000000011111000000000011111000000000000000000000001111111111111111000000000000000001111100000000000000000000000000000000000000000,
354'b000000000000000000000000000000000001111100000000000111111111111100000001111100000000001111100000000011110000000111111110000000111110000000111110000000000000000000000000000000000000111110000000000000000000000111110000000001111000000011110000000000011111000000000000000000000001111111111111111000000000000000001111100000000000000000000000000000000000000000,
354'b000000000000000000000000000000000001111100000000000111111111111100000001111100000000001111100000000011110000000011111100000000111110000000111110000000000000000000000000000000000000111110000000000000000000000111110000000001111100000111110000000000011111000000000000000000000001111100000111111100000000000000001111100000000000000000000000000000000000000000,
354'b000000000000000000000000000000000001111100000000000000000001111100000011111111111111111111110000000011110000000011111100000000111110000000111110000000000000000000000000000000000000011111000000000000000000000111110000000001111100000111110000000000011111000000000000000000000001111100000011111100000000000000001111100000000000000000000000000000000000000000,
354'b000000000000000000000000000000000001111100000000000000000001111100000011111111111111111111110000000011110000000001111100000000111110000000111110000000000000000000000000000000000000011111000000000000000000000111110000000000111100000111100000000000011111000000000000000000000001111100000001111110000000000000001111100000000000000000000000000000000000000000,
354'b000000000000000000000000000000000000111110000000000000000001111100000011111111111111111111110000000011110000000001111000000000111110000000111110000000000000000000000000000000000000011111000000000000000000001111100000000000111110001111100000000000011111000000000000000000000001111100000000111111000000000000001111100000000000000000000000000000000000000000,
354'b000000000000000000000000000000000000111110000000000000000001111100000111111111111111111111111000000011110000000001111000000000111110000000111110000000000000000000000000000000000000011111000000000000000000001111100000000000111110001111100000000000011111000000000000000000000001111100000000011111100000000000001111100000000000000000000000000000000000000000,
354'b000000000000000000000000000000000000111111000000000000000001111100000111110000000000000011111000000011110000000000000000000000111110000000111110000000000000000000000000000000000000001111100000000000000000001111100000000000011110001111000000000000011111000000000000000000000001111100000000001111110000000000000000000000000000000000000000000000000000000000,
354'b000000000000000000000000000000000000011111000000000000000001111100000111100000000000000011111000000011110000000000000000000000111110000000111110000000000000000000000000000000000000001111100000000000000000011111000000000000011111011111000000000000011111000000000000000000000001111100000000001111111000000000000000000000000000000000000000000000000000000000,
354'b000000000000000000000000000000000000011111100000000000000001111100001111100000000000000001111100000011110000000000000000000000111110000000111110000000000000000000000000000000000000001111110000000000000000111111000000000000011111111111000000000000011111000000000000000000000001111100000000000111111000000000000000000000000000000000000000000000000000000000,
354'b000000000000000000000000000000000000001111110000000000000001111100001111100000000000000001111100000011110000000000000000000000111110000000111110000000000000000000000000000000000000000111111000000000000001111110000000000000001111111110000000000000011111000000000000000000000001111100000000000011111100000000000000000000000000000000000000000000000000000000,
354'b000000000000000000000000000000000000001111111000000000000001111100001111000000000000000001111100000011110000000000000000000000111110000000111110000000000000000000000000000000000000000011111100000000000011111110000000000000001111111110000000000000011111000000000000000000000001111100000000000001111110000000000000000000000000000000000000000000000000000000,
354'b000000000000000000000000000000000000000111111110000000000011111100011111000000000000000000111110000011110000000000000000000000111110000000111110000000000000000000000000000000000000000011111111000000000111111100000000000000001111111110000000000000011111000000000000000000000001111100000000000000111111000000001111100000000000000000000000000000000000000000,
354'b000000000000000000000000000000000000000011111111111111111111111100011111000000000000000000111110000011110000000000000000000000111110000000111111111111111111111110000000000000000000000001111111111111111111111000000000000000000111111100000000000000011111111111111111111111000001111100000000000000111111100000001111100000000000000000000000000000000000000000,
354'b000000000000000000000000000000000000000001111111111111111111111100011110000000000000000000111110000011110000000000000000000000111110000000111111111111111111111110000000000000000000000000111111111111111111110000000000000000000111111100000000000000011111111111111111111111000001111100000000000000011111100000001111100000000000000000000000000000000000000000,
354'b000000000000000000000000000000000000000000011111111111111111100000111110000000000000000000011111000011110000000000000000000000111110000000111111111111111111111110000000000000000000000000001111111111111111000000000000000000000111111000000000000000011111111111111111111111000001111100000000000000001111110000001111100000000000000000000000000000000000000000,
354'b000000000000000000000000000000000000000000000111111111111110000000111110000000000000000000011111000011110000000000000000000000111110000000111111111111111111111110000000000000000000000000000011111111111100000000000000000000000011111000000000000000011111111111111111111111000001111100000000000000000111111000001111100000000000000000000000000000000000000000,
354'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000,
354'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000,
354'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000,
354'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000,
354'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000,
354'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000,
354'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000,
354'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000,
354'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000,
354'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000,
354'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000,
354'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000,
354'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000,
354'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000,
354'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000,
354'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000,
354'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000,
354'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000,
354'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000,
354'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000,
354'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000,
354'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000,
354'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000,
354'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000,
354'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000,
354'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000,
354'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000,
354'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000,
354'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000,
354'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000,
354'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000,
354'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000,
354'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000,
354'b111111110000000000011111111000000000000001111111111111110000000011111111000000000001111111100000000000000000001110000000000111100000000001100000000000000000011111111111111111111100000000111111100000000000000000000000111111110000000000000111111111111111100000000111111110000011111111111111111111000000011100000000000011111111000000000011111111111111111111,
354'b111111111111000000011111111111100000000001111111111111110000001111111111111000000111111111111100000000000000001110000000001111100000000011100000000000000000011111111111111111111100000111111111111000000000000000000000111111111111000000000111111111111111100000011111111111110011111111111111111111000000111110000000000011111111111100000011111111111111111111,
354'b111111111111100000011111111111111000000001111111111111110000011111111111111000001111111111111100000000000000001110000000011111000000000111100000000000000000011111111111111111111100001111111111111110000000000000000000111111111111110000000111111111111111100000111111111111110011111111111111111111000000111110000000000011111111111111000011111111111111111111,
354'b111000001111110000011100000011111000000001110000000000000000111110000001111000011111000000111100000000000000001110000000011110000000001111100000000000000000000000000011100000000000011111000000011111000000000000000000111000000111110000000111000000000000000001111100000011110000000000011100000000000001111111000000000011100000011111000000000000011100000000,
354'b111000000011111000011100000000111100000001110000000000000000111100000000011000011110000000001100000000000000001110000000111100000001111111100000000000000000000000000011100000000000111110000000001111000000000000000000111000000001111000000111000000000000000001111000000000110000000000011100000000000001111111000000000011100000000111100000000000011100000000,
354'b111000000001111000011100000000111100000001110000000000000001111000000000000000111100000000000000000000000000001110000001111000000001111111100000000000000000000000000011100000000000111100000000000111100000000000000000111000000001111000000111000000000000000011110000000000000000000000011100000000000001110111000000000011100000000111100000000000011100000000,
354'b111000000000111000011100000000011100000001110000000000000001111000000000000000111100000000000000000000000000001110000011110000000000000011100000000000000000000000000011100000000001111000000000000011100000000000000000111000000000111000000111000000000000000011110000000000000000000000011100000000000011110111100000000011100000000011100000000000011100000000,
354'b111000000000111000011100000000011100000001110000000000000001111000000000000000111100000000000000000000000000001110000111100000000000000011100000000000000000000000000011100000000001111000000000000011110000000000000000111000000000111000000111000000000000000011110000000000000000000000011100000000000011100011100000000011100000000011100000000000011100000000,
354'b111000000000111000011100000000011100000001110000000000000001111000000000000000111100000000000000000000000000001110001111000000000000000011100000000000000000000000000011100000000001110000000000000001110000000000000000111000000000111000000111000000000000000011110000000000000000000000011100000000000011100011100000000011100000000011100000000000011100000000,
354'b111000000000111000011100000000011100000001110000000000000001111100000000000000111110000000000000000000000000001110011110000000000000000011100000000000000000000000000011100000000011110000000000000001110000000000000000111000000000111000000111000000000000000011111000000000000000000000011100000000000111100011110000000011100000000011100000000000011100000000,
354'b111000000000111000011100000000111100000001111111111111110000111110000000000000011111000000000000000000000000001110111100000000000000000011100000000000000000000000000011100000000011110000000000000001111000000000000000111000000001111000000111111111111111000001111100000000000000000000011100000000000111000001110000000011100000000111100000000000011100000000,
354'b111000000001111000011100000001111000000001111111111111110000111111110000000000011111111000000000000000000000001111111000000000000000000011100000000000000000000000000011100000000011110000000000000001111000000000000000111000000011110000000111111111111111000001111111100000000000000000011100000000000111000001110000000011100000001111000000000000011100000000,
354'b111000000011110000011100000011111000000001111111111111110000011111111111000000001111111111100000000000000000001111111100000000000000000011100000000000000000000000000011100000000011110000000000000001111000000000000000111000000111110000000111111111111111000000111111111110000000000000011100000000001111000001111000000011100000011111000000000000011100000000,
354'b111111111111110000011111111111110000000001110000000000000000000111111111110000000011111111111000000000000000001111111100000000000000000011100000000000000000000000000011100000000011110000000000000001111000000000000000111111111111100000000111000000000000000000001111111111100000000000011100000000001110000000111000000011111111111110000000000000011100000000,
354'b111111111111100000011111111111000000000001110000000000000000000000011111111000000000001111111100000000000000001111111110000000000000000011100000000000000000000000000011100000000011110000000000000001111000000000000000111111111110000000000111000000000000000000000000111111110000000000011100000000001110000000111000000011111111111000000000000000011100000000,
354'b111111111110000000011111111111000000000001110000000000000000000000000011111000000000000001111100000000000000001110001111000000000000000011100000000000000000000000000011100000000011110000000000000001111000000000000000111111111110000000000111000000000000000000000000000111110000000000011100000000011110000000111100000011111111111000000000000000011100000000,
354'b111000000000000000011100001111100000000001110000000000000000000000000000111100000000000000011110000000000000001110001111100000000000000011100000000000000000000000000011100000000011110000000000000001111000000000000000111000011111000000000111000000000000000000000000000001111000000000011100000000011111111111111100000011100001111100000000000000011100000000,
354'b111000000000000000011100000111110000000001110000000000000000000000000000111100000000000000011110000000000000001110000111110000000000000011100000000000000000000000000011100000000001110000000000000001110000000000000000111000001111100000000111000000000000000000000000000001111000000000011100000000011111111111111100000011100000111110000000000000011100000000,
354'b111000000000000000011100000011110000000001110000000000000000000000000000011100000000000000001110000000000000001110000011110000000000000011100000000000000000000000000011100000000001111000000000000011110000000000000000111000000111100000000111000000000000000000000000000000111000000000011100000000111111111111111110000011100000011110000000000000011100000000,
354'b111000000000000000011100000001111000000001110000000000000000000000000000011100000000000000001110000000000000001110000001111000000000000011100000000000000000000000000011100000000001111000000000000011110000000000000000111000000011110000000111000000000000000000000000000000111000000000011100000000111000000000001110000011100000001111000000000000011100000000,
354'b111000000000000000011100000000111100000001110000000000000001000000000000111100100000000000011110000000000000001110000001111100000000000011100000000000000000000000000011100000000000111100000000000111100000000000000000111000000001111000000111000000000000000010000000000001111000000000011100000000111000000000001110000011100000000111100000000000011100000000,
354'b111000000000000000011100000000111110000001110000000000000001100000000000111100110000000000011110000000000000001110000000111110000000000011100000000000000000000000000011100000000000111110000000001111100000000000000000111000000001111100000111000000000000000011000000000001111000000000011100000001111000000000001111000011100000000111110000000000011100000000,
354'b111000000000000000011100000000011111000001110000000000000001111000000001111000111100000000111100000000000000001110000000011111000000000011100000000000000000000000000011100000000000011111000000011111000000000000000000111000000000111110000111000000000000000011110000000011110000000000011100000001110000000000000111000011100000000011111000000000011100000000,
354'b111000000000000000011100000000001111000001111111111111110001111111111111110000111111111111111000000000000000001110000000001111000001111111111111000000000000000000000011100000000000001111111111111110000000000000000000111000000000011110000111111111111111100011111111111111100000000000011100000001110000000000000111000011100000000001111000000000011100000000,
354'b111000000000000000011100000000000111100001111111111111110001111111111111100000111111111111110000000000000000001110000000000111100001111111111111000000000000000000000011100000000000000111111111111100000000000000000000111000000000001111000111111111111111100011111111111111000000000000011100000011110000000000000111100011100000000000111100000000011100000000,
354'b111000000000000000011100000000000011110001111111111111110000001111111111000000000111111111100000000000000000001110000000000111110001111111111111000000000000000000000011100000000000000001111111110000000000000000000000111000000000000111100111111111111111100000011111111110000000000000011100000011100000000000000011100011100000000000011110000000011100000000
};


// game over screen message



endmodule
 	
















